
// mux2.v - logic for 2-to-1 multiplexer

module mux2 #(parameter WIDTH = 32) (
    input       [WIDTH-1:0] d0, d1,
    input       sel,
    output      [WIDTH-1:0] y
);

assign y = sel ? d1 : d0;

endmodule

